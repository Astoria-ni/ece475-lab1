//========================================================================
// Lab 1 - Iterative Mul Unit
//========================================================================

`ifndef RISCV_INT_MUL_ITERATIVE_V
`define RISCV_INT_MUL_ITERATIVE_V

module imuldiv_IntMulIterative
(
  input                clk,
  input                reset,

  input  [31:0] mulreq_msg_a,
  input  [31:0] mulreq_msg_b,
  input         mulreq_val,
  output        mulreq_rdy,

  output [63:0] mulresp_msg_result,
  output        mulresp_val,
  input         mulresp_rdy
);

  wire          a_mux_sel;
  wire          b_mux_sel;
  wire          result_mux_sel;
  wire          result_en;
  wire          add_mux_sel;
  wire          cntr_mux_sel;
  wire          sign_en;
  wire          sign_mux_sel;
  wire          b_reg_lsb; //b_reg[0]
  wire    [4:0] counter;

  imuldiv_IntMulIterativeDpath dpath
  (
    .clk                (clk),
    .reset              (reset),
    .mulreq_msg_a       (mulreq_msg_a),
    .mulreq_msg_b       (mulreq_msg_b),
    .mulresp_msg_result (mulresp_msg_result),
    .a_mux_sel          (a_mux_sel),
    .b_mux_sel          (b_mux_sel),
    .result_mux_sel     (result_mux_sel),
    .result_en          (result_en),
    .add_mux_sel        (add_mux_sel),
    .cntr_mux_sel       (cntr_mux_sel),
    .sign_en            (sign_en),
    .sign_mux_sel       (sign_mux_sel),
    .b_reg_lsb          (b_reg_lsb),
    .counter            (counter)
  );

  imuldiv_IntMulIterativeCtrl ctrl
  (
    .clk                (clk),
    .reset              (reset),
    .mulreq_val         (mulreq_val),
    .mulreq_rdy         (mulreq_rdy),
    .mulresp_val        (mulresp_val),
    .mulresp_rdy        (mulresp_rdy),
    .a_mux_sel          (a_mux_sel),
    .b_mux_sel          (b_mux_sel),
    .result_mux_sel     (result_mux_sel),
    .result_en          (result_en),
    .add_mux_sel        (add_mux_sel),
    .cntr_mux_sel       (cntr_mux_sel),
    .sign_en            (sign_en),
    .sign_mux_sel       (sign_mux_sel),
    .b_reg_lsb          (b_reg_lsb),
    .counter            (counter)
  );

endmodule

//------------------------------------------------------------------------
// Datapath
//------------------------------------------------------------------------

module imuldiv_IntMulIterativeDpath
(
  input         clk,
  input         reset,

  input  [31:0] mulreq_msg_a,       // Operand A
  input  [31:0] mulreq_msg_b,       // Operand B
  output [63:0] mulresp_msg_result, // Result of operation

  input         a_mux_sel,
  input         b_mux_sel,
  input         result_mux_sel,
  input         result_en,
  input         add_mux_sel,
  input         cntr_mux_sel,
  input         sign_en,
  input         sign_mux_sel,

  output        b_reg_lsb,
  output  [4:0] counter
);

  assign mulresp_msg_result = 64'b0;
  assign b_reg_lsb          = 1'b0;
  assign counter            = 5'b0;
  /*
  //----------------------------------------------------------------------
  // Sequential Logic
  //----------------------------------------------------------------------

  reg  [63:0] a_reg;       // Register for storing operand A
  reg  [31:0] b_reg;       // Register for storing operand B
  reg         val_reg;     // Register for storing valid bit

  always @( posedge clk ) begin

    // Stall the pipeline if the response interface is not ready
    if ( mulresp_rdy ) begin
      a_reg   <= mulreq_msg_a;
      b_reg   <= mulreq_msg_b;
      val_reg <= mulreq_val;
    end

  end

  //----------------------------------------------------------------------
  // Combinational Logic
  //----------------------------------------------------------------------

  // Extract sign bits

  wire sign_bit_a = a_reg[31];
  wire sign_bit_b = b_reg[31];

  // Unsign operands if necessary

  wire [31:0] unsigned_a = ( sign_bit_a ) ? (~a_reg + 1'b1) : a_reg;
  wire [31:0] unsigned_b = ( sign_bit_b ) ? (~b_reg + 1'b1) : b_reg;

  // Computation logic

  wire [63:0] unsigned_result = unsigned_a * unsigned_b;

  // Determine whether or not result is signed. Usually the result is
  // signed if one and only one of the input operands is signed. In other
  // words, the result is signed if the xor of the sign bits of the input
  // operands is true. Remainder opeartions are a bit trickier, and here
  // we simply assume that the result is signed if the dividend for the
  // rem operation is signed.

  wire is_result_signed = sign_bit_a ^ sign_bit_b;

  assign mulresp_msg_result
    = ( is_result_signed ) ? (~unsigned_result + 1'b1) : unsigned_result;

  // Set the val/rdy signals. The request is ready when the response is
  // ready, and the response is valid when there is valid data in the
  // input registers.

  assign mulreq_rdy  = mulresp_rdy;
  assign mulresp_val = val_reg;
  */
endmodule

//------------------------------------------------------------------------
// Control Logic
//------------------------------------------------------------------------

module imuldiv_IntMulIterativeCtrl
(
  input         clk,
  input         reset,

  input         mulreq_val,
  output        mulreq_rdy,
  output        mulresp_val,
  input         mulresp_rdy,

  output        a_mux_sel,
  output        b_mux_sel,
  output        result_mux_sel,
  output        result_en,
  output        add_mux_sel,
  output        cntr_mux_sel,
  output        sign_en,
  output        sign_mux_sel,

  input         b_reg_lsb,
  input   [4:0] counter
);
  
  assign mulreq_rdy = 1'b1;
  assign mulresp_val= 1'b0;

  assign a_mux_sel  = 1'b0;
  assign b_mux_sel  = 1'b0;
  assign result_mux_sel = 1'b0;
  assign result_en  = 1'b0;
  assign add_mux_sel = 1'b0;
  assign cntr_mux_sel = 1'b0;
  assign sign_en     = 1'b0;
  assign sign_mux_sel = 1'b0;

endmodule

`endif
